library verilog;
use verilog.vl_types.all;
entity proyecto1_vlg_vec_tst is
end proyecto1_vlg_vec_tst;
